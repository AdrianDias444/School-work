* ============================================
* 1. FUNCIONAMENTO BÁSICO DO RETIFICADOR
*    (Onda completa com center-tap)
* ============================================
* Objetivo: Validar o princípio de funcionamento
* Saída formatada para gnuplot
* ============================================

* 1.1 FONTES DE ENTRADA
Vin entrada 0 SIN(0 10 60)                   ; Fonte primária: 10Vp, 60Hz
B1 sec1 0 V = +5*sin(2*3.14159*60*time)     ; Secundário 1: +5V (center-tap)
B2 sec2 0 V = -5*sin(2*3.14159*60*time)     ; Secundário 2: -5V (180° defasado)

* 1.2 RETIFICADOR DE ONDA COMPLETA
D1 sec1 saida 1N4007                        ; Diodo superior
D2 sec2 saida 1N4007                        ; Diodo inferior
.model 1N4007 D(IS=14.11e-9 N=1.984 RS=0.1) ; Modelo real do diodo

* 1.3 CARGA
R_carga saida 0 1k                          ; Resistência de carga

* ============================================
* 2. ANÁLISE TRANSIENTE
* ============================================
.tran 0.1ms 100ms                           ; 100ms (~6 ciclos de 60Hz)

* ============================================
* 3. MEDIÇÕES (opcional, para relatório)
* ============================================
.measure tran Vdc_medio avg V(saida) from=50ms to=100ms
.measure tran Vripple_pp pp V(saida) from=50ms to=100ms
.measure tran freq_ripple param 120         ; Teórico: 2×60Hz = 120Hz

* ============================================
* 4. SAÍDA PARA GNUPLOT
* ============================================
* Opção para manter todos os pontos
.option plotwinsize=0

* Salvar dados em formato tabular
.print tran v(entrada) v(saida)
* Ou, alternativamente, salvar em arquivo específico:
* .write dados_retificador.dat v(entrada) v(saida)

* ============================================
* 5. FIM DA NETLIST
* ============================================
.end
