* ============================================
* 3. FILTRO CAPACITIVO
* ============================================
* Objetivo: Reduzir ripple com capacitor

Vin entrada 0 SIN(0 10 60)
B1 sec1 0 V = +5*sin(2*3.14159*60*time)
B2 sec2 0 V = -5*sin(2*3.14159*60*time)
D1 sec1 saida 1N4007
D2 sec2 saida 1N4007
.model 1N4007 D(IS=14.11e-9 N=1.984 RS=0.1)
R_carga saida 0 1k

* CAPACITOR DE FILTRO (alterar manualmente para cada teste)
C_filtro saida 0 100u  ; TESTAR: 10u, 100u, 1000u

.tran 0.1ms 100ms

.measure tran Vdc avg V(saida) from=50ms to=100ms
.measure tran Vripple pp V(saida) from=50ms to=100ms
.measure tran Idiodo_pico max I(D1) from=0 to=100ms

.print tran Vdc Vripple Idiodo_pico
.plot tran v(saida)

.end
