* FALHA: DIODO D1 ABERTO
Vin entrada 0 SIN(0 10 60)
B1 sec1 0 V = +5*sin(2*3.14159*60*time)
B2 sec2 0 V = -5*sin(2*3.14159*60*time)

* APENAS D2 FUNCIONA - D1 ESTÁ ABERTO
D2 sec2 saida 1N4007    ; Apenas este diodo

.model 1N4007 D(IS=14.11e-9 N=1.984 RS=0.1)
R_carga saida 0 1k
C_filtro saida 0 100u

.tran 0.1ms 100ms

.measure tran Vdc_falha avg V(saida) from=50ms to=100ms
.measure tran Vripple_falha pp V(saida) from=50ms to=100ms

.print tran Vdc_falha Vripple_falha
.plot tran v(saida)

.end
